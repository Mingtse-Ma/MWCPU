//总线顶层模块
module（）；
endmodule